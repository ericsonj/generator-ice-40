/**
 * File:   <%= projectName %>.v
 * Author: <%= username %>
 * Email:  <%= email %>
 * 
 * Created on <%= datetime %>
 */

module <%= projectName %> (/*PORTS*/);
endmodule // <%= projectName %>
